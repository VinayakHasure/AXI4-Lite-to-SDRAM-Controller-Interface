`include "uvm_macros.svh"
import uvm_pkg::*;

`include "../AXI/AXI_Interface.sv"
`include "../AXI/AXI_Packet.sv"
`include "../AXI/AXI_Base_Sequence.sv"
`include "../AXI/AXI_Sequence.sv"
`include "../AXI/AXI_Sequencer.sv"
`include "../AXI/AXI_Driver.sv"
`include "../AXI/AXI_Monitor.sv"
`include "../AXI/AXI_Agent.sv"
`include "../SDRAM/SDRAM_Interface.sv"
`include "../SDRAM/SDRAM_Packet.sv"
`include "../SDRAM/SDRAM_base_Sequence.sv"
`include "../SDRAM/SDRAM_Sequence.sv"
`include "../SDRAM/SDRAM_Sequencer.sv"
`include "../SDRAM/SDRAM_Driver.sv"
`include "../SDRAM/SDRAM_Monitor.sv"
`include "../SDRAM/SDRAM_Agent.sv"
`include "AXI_SDRAM_Scoreboard.sv"
`include "AXI_SDRAM_Coverage.sv"
`include "AXI2SDRAM_Environment.sv"
`include "AXI_SDRAM_Test.sv"
// `include "../../Design/AXI2SDRAM_Wrapper/async_fifo.sv"
// `include "../../Design/AXI2SDRAM_Wrapper/axi_slave_fsm.sv"
// `include "../../Design/AXI2SDRAM_Wrapper/fifo.sv"
// `include "../../Design/AXI2SDRAM_Wrapper/SDRAM_Controller.sv"
// `include "../../Design/AXI2SDRAM_Wrapper/axi2sdram_wrapper.sv"
// `include "../../Design/sdram_sim_model/mt48lc16m16a2.v"
